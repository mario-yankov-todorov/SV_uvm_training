module memory_driver
    (
      input clk,
      input rst,
      input data_in,
      output full
    );

endmodule
