interface dut_if;
  
   logic   clk        ;
   logic   rst        ;
   logic   button     ;
   
   logic   MEM_FULL   ;
   
endinterface