// When the test bench is fully developed here will be the design of the memory_driver
module memory_driver 
  (
      dut_if   dif   ;
  );
  
  
endmodule