module assertion_penable
   (
       input   clk          ,
       input   PWRITE       ,
       input   PSEL         ,
       input   PENABLE            
   );
  
  
endmodule